module local_branch_predictor #
(
    parameter ADDR_WIDTH = 32
)
(
    input wire clk,
    input wire sel,
    
);
    
endmodule
