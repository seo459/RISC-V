module branch_top #
(
    parameter ADDR_WIDTH = 32
)
(
    input wire clk,
    input wire sel,
    
);
    
endmodule
